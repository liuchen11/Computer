library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity VGA is
   Port (
		clk	: in	std_logic;
      rst	: in	std_logic;
      R		: out	std_logic_vector(2 downto 0);
      G		: out	std_logic_vector(2 downto 0);
      B		: out	std_logic_vector(2 downto 0);
      Hs		: out	std_logic;
      Vs		: out	std_logic
	);
end VGA;
architecture Behavioral of VGA is
signal stdclk	:std_logic:='0';
signal div		:std_logic:='0';
shared variable col:integer range 0 to 800:=0;
shared variable row:integer range 0 to 525:=0;

begin
divide:process(clk)
begin
	if rising_edge(clk) then
		stdclk<=not stdclk;
	end if;
end process;
scan:process(stdclk,rst)
begin
	if rst='0' then
		col:=0;
		row:=0;
	elsif rising_edge(stdclk) then
		case row is		
			when 180=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 181=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 182=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 183=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 184=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 185=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 186=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 187=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 188=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 189=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 190=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 191=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 192=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 193=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 194=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "010";G <= "010";B <= "011";
					when 252=>
						R <= "111";G <= "111";B <= "111";
					when 253=>
						R <= "111";G <= "111";B <= "111";
					when 254=>
						R <= "111";G <= "111";B <= "111";
					when 255=>
						R <= "111";G <= "111";B <= "111";
					when 256=>
						R <= "111";G <= "111";B <= "111";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "111";
					when 259=>
						R <= "111";G <= "111";B <= "111";
					when 260=>
						R <= "111";G <= "111";B <= "111";
					when 261=>
						R <= "111";G <= "111";B <= "111";
					when 262=>
						R <= "111";G <= "111";B <= "111";
					when 263=>
						R <= "111";G <= "111";B <= "111";
					when 264=>
						R <= "100";G <= "011";B <= "010";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "101";B <= "100";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "001";G <= "010";B <= "011";
					when 285=>
						R <= "111";G <= "111";B <= "111";
					when 286=>
						R <= "111";G <= "111";B <= "111";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "111";G <= "111";B <= "111";
					when 289=>
						R <= "111";G <= "111";B <= "111";
					when 290=>
						R <= "101";G <= "100";B <= "011";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "111";B <= "111";
					when 296=>
						R <= "110";G <= "110";B <= "101";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "101";G <= "110";B <= "110";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "101";B <= "100";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "101";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "111";B <= "111";
					when 316=>
						R <= "111";G <= "111";B <= "111";
					when 317=>
						R <= "111";G <= "111";B <= "111";
					when 318=>
						R <= "111";G <= "111";B <= "111";
					when 319=>
						R <= "111";G <= "111";B <= "111";
					when 320=>
						R <= "111";G <= "111";B <= "111";
					when 321=>
						R <= "111";G <= "110";B <= "110";
					when 322=>
						R <= "001";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "001";
					when 333=>
						R <= "110";G <= "111";B <= "111";
					when 334=>
						R <= "111";G <= "111";B <= "111";
					when 335=>
						R <= "111";G <= "111";B <= "111";
					when 336=>
						R <= "001";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "111";G <= "111";B <= "111";
					when 348=>
						R <= "111";G <= "111";B <= "111";
					when 349=>
						R <= "111";G <= "111";B <= "111";
					when 350=>
						R <= "111";G <= "111";B <= "111";
					when 351=>
						R <= "111";G <= "111";B <= "111";
					when 352=>
						R <= "111";G <= "111";B <= "111";
					when 353=>
						R <= "111";G <= "111";B <= "111";
					when 354=>
						R <= "001";G <= "001";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 195=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "010";G <= "010";B <= "010";
					when 252=>
						R <= "111";G <= "111";B <= "111";
					when 253=>
						R <= "111";G <= "111";B <= "111";
					when 254=>
						R <= "111";G <= "111";B <= "111";
					when 255=>
						R <= "111";G <= "111";B <= "111";
					when 256=>
						R <= "111";G <= "111";B <= "111";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "111";
					when 259=>
						R <= "111";G <= "111";B <= "111";
					when 260=>
						R <= "111";G <= "111";B <= "111";
					when 261=>
						R <= "111";G <= "111";B <= "111";
					when 262=>
						R <= "111";G <= "111";B <= "111";
					when 263=>
						R <= "111";G <= "111";B <= "111";
					when 264=>
						R <= "100";G <= "011";B <= "010";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "101";
					when 270=>
						R <= "001";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "010";G <= "010";B <= "011";
					when 285=>
						R <= "111";G <= "111";B <= "111";
					when 286=>
						R <= "111";G <= "111";B <= "111";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "111";G <= "111";B <= "111";
					when 289=>
						R <= "111";G <= "111";B <= "111";
					when 290=>
						R <= "101";G <= "100";B <= "100";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "111";B <= "111";
					when 296=>
						R <= "111";G <= "111";B <= "111";
					when 297=>
						R <= "100";G <= "011";B <= "010";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "001";
					when 306=>
						R <= "101";G <= "110";B <= "110";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "011";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "101";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "111";B <= "111";
					when 316=>
						R <= "111";G <= "111";B <= "111";
					when 317=>
						R <= "111";G <= "111";B <= "111";
					when 318=>
						R <= "111";G <= "111";B <= "111";
					when 319=>
						R <= "111";G <= "111";B <= "111";
					when 320=>
						R <= "111";G <= "111";B <= "111";
					when 321=>
						R <= "111";G <= "111";B <= "111";
					when 322=>
						R <= "111";G <= "111";B <= "111";
					when 323=>
						R <= "101";G <= "100";B <= "100";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "001";G <= "010";B <= "011";
					when 333=>
						R <= "111";G <= "111";B <= "111";
					when 334=>
						R <= "111";G <= "111";B <= "111";
					when 335=>
						R <= "111";G <= "111";B <= "111";
					when 336=>
						R <= "100";G <= "011";B <= "010";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "100";G <= "101";B <= "110";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "111";G <= "111";B <= "111";
					when 348=>
						R <= "111";G <= "111";B <= "111";
					when 349=>
						R <= "111";G <= "111";B <= "111";
					when 350=>
						R <= "111";G <= "111";B <= "111";
					when 351=>
						R <= "111";G <= "111";B <= "111";
					when 352=>
						R <= "111";G <= "111";B <= "111";
					when 353=>
						R <= "111";G <= "111";B <= "111";
					when 354=>
						R <= "111";G <= "111";B <= "111";
					when 355=>
						R <= "111";G <= "111";B <= "111";
					when 356=>
						R <= "010";G <= "010";B <= "010";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 196=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "001";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "111";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "101";
					when 270=>
						R <= "001";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "110";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "001";
					when 293=>
						R <= "011";G <= "100";B <= "101";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "111";B <= "111";
					when 296=>
						R <= "111";G <= "111";B <= "111";
					when 297=>
						R <= "111";G <= "111";B <= "110";
					when 298=>
						R <= "001";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "001";
					when 306=>
						R <= "101";G <= "110";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "100";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "101";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "001";G <= "001";B <= "010";
					when 321=>
						R <= "111";G <= "111";B <= "111";
					when 322=>
						R <= "111";G <= "111";B <= "111";
					when 323=>
						R <= "111";G <= "111";B <= "111";
					when 324=>
						R <= "010";G <= "010";B <= "001";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "100";G <= "101";B <= "101";
					when 333=>
						R <= "111";G <= "111";B <= "111";
					when 334=>
						R <= "110";G <= "110";B <= "111";
					when 335=>
						R <= "111";G <= "111";B <= "111";
					when 336=>
						R <= "110";G <= "110";B <= "101";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "110";B <= "101";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "011";G <= "100";B <= "100";
					when 354=>
						R <= "111";G <= "111";B <= "111";
					when 355=>
						R <= "111";G <= "111";B <= "111";
					when 356=>
						R <= "111";G <= "111";B <= "111";
					when 357=>
						R <= "100";G <= "011";B <= "010";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 197=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "001";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "110";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "001";
					when 293=>
						R <= "011";G <= "100";B <= "101";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "111";B <= "111";
					when 296=>
						R <= "111";G <= "111";B <= "111";
					when 297=>
						R <= "111";G <= "111";B <= "111";
					when 298=>
						R <= "110";G <= "101";B <= "101";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "001";
					when 306=>
						R <= "101";G <= "110";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "100";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "111";B <= "110";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "001";
					when 322=>
						R <= "110";G <= "111";B <= "111";
					when 323=>
						R <= "111";G <= "111";B <= "111";
					when 324=>
						R <= "110";G <= "101";B <= "101";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "001";G <= "001";B <= "010";
					when 332=>
						R <= "111";G <= "111";B <= "111";
					when 333=>
						R <= "111";G <= "111";B <= "111";
					when 334=>
						R <= "010";G <= "010";B <= "011";
					when 335=>
						R <= "111";G <= "111";B <= "111";
					when 336=>
						R <= "111";G <= "111";B <= "110";
					when 337=>
						R <= "011";G <= "010";B <= "001";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "001";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "110";B <= "100";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "001";
					when 355=>
						R <= "101";G <= "110";B <= "110";
					when 356=>
						R <= "111";G <= "111";B <= "111";
					when 357=>
						R <= "111";G <= "111";B <= "111";
					when 358=>
						R <= "100";G <= "011";B <= "010";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 198=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "001";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "110";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "001";
					when 293=>
						R <= "011";G <= "100";B <= "101";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "110";
					when 296=>
						R <= "011";G <= "011";B <= "011";
					when 297=>
						R <= "111";G <= "111";B <= "111";
					when 298=>
						R <= "111";G <= "111";B <= "111";
					when 299=>
						R <= "100";G <= "011";B <= "010";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "101";G <= "110";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "100";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "101";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "100";G <= "101";B <= "110";
					when 323=>
						R <= "111";G <= "111";B <= "111";
					when 324=>
						R <= "111";G <= "110";B <= "110";
					when 325=>
						R <= "001";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "011";G <= "100";B <= "100";
					when 332=>
						R <= "111";G <= "111";B <= "111";
					when 333=>
						R <= "110";G <= "110";B <= "101";
					when 334=>
						R <= "000";G <= "000";B <= "001";
					when 335=>
						R <= "101";G <= "110";B <= "111";
					when 336=>
						R <= "111";G <= "111";B <= "111";
					when 337=>
						R <= "101";G <= "101";B <= "100";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "001";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "110";B <= "101";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "101";G <= "110";B <= "110";
					when 357=>
						R <= "111";G <= "111";B <= "111";
					when 358=>
						R <= "111";G <= "111";B <= "111";
					when 359=>
						R <= "001";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 199=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "101";
					when 270=>
						R <= "001";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "110";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "001";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "110";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "101";G <= "101";B <= "101";
					when 298=>
						R <= "111";G <= "111";B <= "111";
					when 299=>
						R <= "111";G <= "111";B <= "111";
					when 300=>
						R <= "001";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "101";G <= "110";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "100";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "110";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "011";G <= "100";B <= "100";
					when 323=>
						R <= "111";G <= "111";B <= "111";
					when 324=>
						R <= "111";G <= "111";B <= "110";
					when 325=>
						R <= "001";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "001";
					when 331=>
						R <= "101";G <= "110";B <= "110";
					when 332=>
						R <= "111";G <= "111";B <= "111";
					when 333=>
						R <= "100";G <= "011";B <= "010";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "011";G <= "100";B <= "101";
					when 336=>
						R <= "111";G <= "111";B <= "111";
					when 337=>
						R <= "111";G <= "110";B <= "110";
					when 338=>
						R <= "001";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "001";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "101";B <= "101";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "001";B <= "010";
					when 357=>
						R <= "110";G <= "111";B <= "111";
					when 358=>
						R <= "111";G <= "111";B <= "111";
					when 359=>
						R <= "101";G <= "100";B <= "011";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 200=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "001";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "110";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "110";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "110";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "001";
					when 298=>
						R <= "110";G <= "111";B <= "111";
					when 299=>
						R <= "111";G <= "111";B <= "111";
					when 300=>
						R <= "110";G <= "101";B <= "101";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "101";G <= "110";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "100";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "101";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "100";G <= "101";B <= "101";
					when 323=>
						R <= "111";G <= "111";B <= "111";
					when 324=>
						R <= "111";G <= "110";B <= "101";
					when 325=>
						R <= "001";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "001";G <= "010";B <= "011";
					when 331=>
						R <= "111";G <= "111";B <= "111";
					when 332=>
						R <= "111";G <= "111";B <= "110";
					when 333=>
						R <= "001";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "001";G <= "001";B <= "010";
					when 336=>
						R <= "111";G <= "111";B <= "111";
					when 337=>
						R <= "111";G <= "111";B <= "111";
					when 338=>
						R <= "100";G <= "011";B <= "010";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "001";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "101";B <= "101";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "001";
					when 357=>
						R <= "101";G <= "110";B <= "111";
					when 358=>
						R <= "111";G <= "111";B <= "110";
					when 359=>
						R <= "110";G <= "110";B <= "100";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 201=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "110";G <= "110";B <= "110";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "110";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "110";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "001";G <= "010";B <= "011";
					when 299=>
						R <= "111";G <= "111";B <= "111";
					when 300=>
						R <= "111";G <= "111";B <= "111";
					when 301=>
						R <= "100";G <= "011";B <= "010";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "101";G <= "110";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "100";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "110";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "001";G <= "001";B <= "010";
					when 322=>
						R <= "111";G <= "111";B <= "111";
					when 323=>
						R <= "111";G <= "111";B <= "111";
					when 324=>
						R <= "101";G <= "100";B <= "100";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "100";G <= "101";B <= "101";
					when 331=>
						R <= "111";G <= "111";B <= "111";
					when 332=>
						R <= "110";G <= "110";B <= "101";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "001";
					when 336=>
						R <= "101";G <= "110";B <= "111";
					when 337=>
						R <= "111";G <= "111";B <= "111";
					when 338=>
						R <= "110";G <= "110";B <= "101";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "001";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "101";B <= "101";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "001";
					when 357=>
						R <= "100";G <= "101";B <= "110";
					when 358=>
						R <= "111";G <= "111";B <= "111";
					when 359=>
						R <= "111";G <= "110";B <= "101";
					when 360=>
						R <= "001";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 202=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "111";B <= "110";
					when 270=>
						R <= "111";G <= "111";B <= "111";
					when 271=>
						R <= "111";G <= "111";B <= "111";
					when 272=>
						R <= "111";G <= "111";B <= "111";
					when 273=>
						R <= "111";G <= "111";B <= "111";
					when 274=>
						R <= "111";G <= "111";B <= "111";
					when 275=>
						R <= "111";G <= "111";B <= "111";
					when 276=>
						R <= "111";G <= "111";B <= "111";
					when 277=>
						R <= "111";G <= "111";B <= "111";
					when 278=>
						R <= "111";G <= "111";B <= "111";
					when 279=>
						R <= "111";G <= "111";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "110";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "110";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "110";
					when 296=>
						R <= "001";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "001";
					when 299=>
						R <= "100";G <= "101";B <= "110";
					when 300=>
						R <= "111";G <= "111";B <= "111";
					when 301=>
						R <= "111";G <= "111";B <= "111";
					when 302=>
						R <= "001";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "001";
					when 306=>
						R <= "101";G <= "110";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "011";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "110";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "001";G <= "010";B <= "010";
					when 321=>
						R <= "111";G <= "111";B <= "111";
					when 322=>
						R <= "111";G <= "111";B <= "111";
					when 323=>
						R <= "111";G <= "111";B <= "111";
					when 324=>
						R <= "001";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "001";
					when 330=>
						R <= "110";G <= "111";B <= "111";
					when 331=>
						R <= "111";G <= "111";B <= "111";
					when 332=>
						R <= "100";G <= "011";B <= "010";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "001";G <= "010";B <= "011";
					when 337=>
						R <= "111";G <= "111";B <= "111";
					when 338=>
						R <= "111";G <= "111";B <= "110";
					when 339=>
						R <= "001";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "001";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "101";B <= "100";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "001";
					when 357=>
						R <= "011";G <= "100";B <= "100";
					when 358=>
						R <= "111";G <= "111";B <= "111";
					when 359=>
						R <= "111";G <= "111";B <= "110";
					when 360=>
						R <= "001";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 203=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "111";B <= "111";
					when 270=>
						R <= "111";G <= "111";B <= "111";
					when 271=>
						R <= "111";G <= "111";B <= "111";
					when 272=>
						R <= "111";G <= "111";B <= "111";
					when 273=>
						R <= "111";G <= "111";B <= "111";
					when 274=>
						R <= "111";G <= "111";B <= "111";
					when 275=>
						R <= "111";G <= "111";B <= "111";
					when 276=>
						R <= "111";G <= "111";B <= "111";
					when 277=>
						R <= "111";G <= "111";B <= "111";
					when 278=>
						R <= "111";G <= "111";B <= "111";
					when 279=>
						R <= "111";G <= "111";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "110";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "101";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "001";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "110";
					when 296=>
						R <= "001";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "001";
					when 300=>
						R <= "110";G <= "111";B <= "111";
					when 301=>
						R <= "111";G <= "111";B <= "111";
					when 302=>
						R <= "110";G <= "101";B <= "101";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "001";
					when 306=>
						R <= "101";G <= "110";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "011";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "111";B <= "111";
					when 316=>
						R <= "111";G <= "111";B <= "111";
					when 317=>
						R <= "111";G <= "111";B <= "111";
					when 318=>
						R <= "111";G <= "111";B <= "111";
					when 319=>
						R <= "111";G <= "111";B <= "111";
					when 320=>
						R <= "111";G <= "111";B <= "111";
					when 321=>
						R <= "111";G <= "111";B <= "111";
					when 322=>
						R <= "111";G <= "111";B <= "111";
					when 323=>
						R <= "001";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "001";
					when 329=>
						R <= "011";G <= "100";B <= "100";
					when 330=>
						R <= "111";G <= "111";B <= "111";
					when 331=>
						R <= "111";G <= "111";B <= "111";
					when 332=>
						R <= "001";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "001";
					when 337=>
						R <= "110";G <= "111";B <= "111";
					when 338=>
						R <= "111";G <= "111";B <= "111";
					when 339=>
						R <= "101";G <= "100";B <= "011";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "001";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "101";B <= "100";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "001";
					when 357=>
						R <= "011";G <= "100";B <= "100";
					when 358=>
						R <= "111";G <= "111";B <= "111";
					when 359=>
						R <= "111";G <= "111";B <= "110";
					when 360=>
						R <= "001";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 204=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "110";G <= "110";B <= "110";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "101";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "001";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "110";
					when 296=>
						R <= "001";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "001";G <= "010";B <= "011";
					when 301=>
						R <= "111";G <= "111";B <= "111";
					when 302=>
						R <= "111";G <= "111";B <= "111";
					when 303=>
						R <= "100";G <= "011";B <= "010";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "101";G <= "110";B <= "110";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "011";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "111";B <= "111";
					when 316=>
						R <= "111";G <= "111";B <= "111";
					when 317=>
						R <= "111";G <= "111";B <= "111";
					when 318=>
						R <= "111";G <= "111";B <= "111";
					when 319=>
						R <= "111";G <= "111";B <= "111";
					when 320=>
						R <= "111";G <= "111";B <= "111";
					when 321=>
						R <= "011";G <= "011";B <= "010";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "001";
					when 329=>
						R <= "101";G <= "110";B <= "111";
					when 330=>
						R <= "111";G <= "111";B <= "111";
					when 331=>
						R <= "101";G <= "100";B <= "100";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "100";G <= "101";B <= "101";
					when 338=>
						R <= "111";G <= "111";B <= "111";
					when 339=>
						R <= "111";G <= "110";B <= "110";
					when 340=>
						R <= "001";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "001";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "111";G <= "110";B <= "101";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "001";
					when 357=>
						R <= "100";G <= "101";B <= "110";
					when 358=>
						R <= "111";G <= "111";B <= "111";
					when 359=>
						R <= "111";G <= "110";B <= "101";
					when 360=>
						R <= "001";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 205=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "101";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "001";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "101";
					when 296=>
						R <= "001";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "100";G <= "101";B <= "101";
					when 302=>
						R <= "111";G <= "111";B <= "111";
					when 303=>
						R <= "111";G <= "111";B <= "111";
					when 304=>
						R <= "001";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "101";G <= "110";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "011";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "110";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "001";B <= "010";
					when 329=>
						R <= "110";G <= "111";B <= "111";
					when 330=>
						R <= "111";G <= "111";B <= "111";
					when 331=>
						R <= "111";G <= "111";B <= "111";
					when 332=>
						R <= "111";G <= "111";B <= "111";
					when 333=>
						R <= "111";G <= "111";B <= "111";
					when 334=>
						R <= "111";G <= "111";B <= "111";
					when 335=>
						R <= "111";G <= "111";B <= "111";
					when 336=>
						R <= "111";G <= "111";B <= "111";
					when 337=>
						R <= "111";G <= "111";B <= "111";
					when 338=>
						R <= "111";G <= "111";B <= "111";
					when 339=>
						R <= "111";G <= "111";B <= "111";
					when 340=>
						R <= "011";G <= "010";B <= "001";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "001";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "110";B <= "101";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "001";
					when 357=>
						R <= "101";G <= "110";B <= "111";
					when 358=>
						R <= "111";G <= "111";B <= "111";
					when 359=>
						R <= "110";G <= "101";B <= "100";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 206=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "110";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "001";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "101";
					when 296=>
						R <= "001";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "110";G <= "111";B <= "111";
					when 303=>
						R <= "111";G <= "111";B <= "111";
					when 304=>
						R <= "110";G <= "110";B <= "101";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "100";G <= "101";B <= "101";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "100";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "110";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "100";G <= "101";B <= "110";
					when 329=>
						R <= "111";G <= "111";B <= "111";
					when 330=>
						R <= "111";G <= "111";B <= "111";
					when 331=>
						R <= "111";G <= "111";B <= "111";
					when 332=>
						R <= "111";G <= "111";B <= "111";
					when 333=>
						R <= "111";G <= "111";B <= "111";
					when 334=>
						R <= "111";G <= "111";B <= "111";
					when 335=>
						R <= "111";G <= "111";B <= "111";
					when 336=>
						R <= "111";G <= "111";B <= "111";
					when 337=>
						R <= "111";G <= "111";B <= "111";
					when 338=>
						R <= "111";G <= "111";B <= "111";
					when 339=>
						R <= "111";G <= "111";B <= "111";
					when 340=>
						R <= "110";G <= "101";B <= "101";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "110";B <= "101";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "001";G <= "010";B <= "011";
					when 357=>
						R <= "111";G <= "111";B <= "111";
					when 358=>
						R <= "111";G <= "111";B <= "110";
					when 359=>
						R <= "100";G <= "011";B <= "010";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 207=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "001";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "101";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "001";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "110";
					when 296=>
						R <= "001";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "010";G <= "010";B <= "011";
					when 303=>
						R <= "111";G <= "111";B <= "111";
					when 304=>
						R <= "111";G <= "111";B <= "111";
					when 305=>
						R <= "011";G <= "011";B <= "011";
					when 306=>
						R <= "101";G <= "101";B <= "101";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "100";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "101";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "001";
					when 328=>
						R <= "110";G <= "111";B <= "111";
					when 329=>
						R <= "111";G <= "111";B <= "111";
					when 330=>
						R <= "101";G <= "100";B <= "100";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "011";G <= "100";B <= "100";
					when 339=>
						R <= "111";G <= "111";B <= "111";
					when 340=>
						R <= "111";G <= "111";B <= "111";
					when 341=>
						R <= "001";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "101";B <= "100";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "101";G <= "110";B <= "110";
					when 357=>
						R <= "111";G <= "111";B <= "111";
					when 358=>
						R <= "111";G <= "110";B <= "110";
					when 359=>
						R <= "001";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 208=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "001";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "110";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "110";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "101";
					when 296=>
						R <= "001";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "011";G <= "100";B <= "100";
					when 304=>
						R <= "111";G <= "111";B <= "111";
					when 305=>
						R <= "111";G <= "111";B <= "111";
					when 306=>
						R <= "101";G <= "101";B <= "110";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "011";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "101";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "001";
					when 327=>
						R <= "001";G <= "010";B <= "011";
					when 328=>
						R <= "111";G <= "111";B <= "111";
					when 329=>
						R <= "111";G <= "111";B <= "111";
					when 330=>
						R <= "011";G <= "010";B <= "001";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "001";B <= "010";
					when 339=>
						R <= "111";G <= "111";B <= "111";
					when 340=>
						R <= "111";G <= "111";B <= "111";
					when 341=>
						R <= "100";G <= "011";B <= "010";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "110";B <= "101";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "110";G <= "110";B <= "110";
					when 356=>
						R <= "111";G <= "111";B <= "111";
					when 357=>
						R <= "111";G <= "111";B <= "111";
					when 358=>
						R <= "010";G <= "010";B <= "001";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 209=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "001";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "100";G <= "101";B <= "110";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "110";G <= "110";B <= "101";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "110";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "001";
					when 304=>
						R <= "101";G <= "110";B <= "110";
					when 305=>
						R <= "111";G <= "111";B <= "111";
					when 306=>
						R <= "111";G <= "111";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "011";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "101";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "001";
					when 327=>
						R <= "101";G <= "110";B <= "111";
					when 328=>
						R <= "111";G <= "111";B <= "111";
					when 329=>
						R <= "111";G <= "110";B <= "101";
					when 330=>
						R <= "001";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "001";
					when 339=>
						R <= "101";G <= "110";B <= "111";
					when 340=>
						R <= "111";G <= "111";B <= "111";
					when 341=>
						R <= "111";G <= "110";B <= "110";
					when 342=>
						R <= "001";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "100";G <= "101";B <= "101";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "110";B <= "101";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "100";G <= "101";B <= "101";
					when 354=>
						R <= "111";G <= "111";B <= "111";
					when 355=>
						R <= "111";G <= "111";B <= "111";
					when 356=>
						R <= "111";G <= "111";B <= "111";
					when 357=>
						R <= "010";G <= "010";B <= "001";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "001";G <= "001";B <= "010";
					when 363=>
						R <= "111";G <= "111";B <= "111";
					when 364=>
						R <= "111";G <= "111";B <= "111";
					when 365=>
						R <= "011";G <= "010";B <= "001";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "001";B <= "010";
					when 369=>
						R <= "111";G <= "111";B <= "111";
					when 370=>
						R <= "111";G <= "111";B <= "111";
					when 371=>
						R <= "010";G <= "010";B <= "001";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "001";B <= "010";
					when 375=>
						R <= "111";G <= "111";B <= "111";
					when 376=>
						R <= "111";G <= "111";B <= "111";
					when 377=>
						R <= "010";G <= "010";B <= "001";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 210=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "110";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "001";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "101";
					when 270=>
						R <= "001";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "001";
					when 279=>
						R <= "101";G <= "110";B <= "111";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "011";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "001";G <= "010";B <= "011";
					when 285=>
						R <= "111";G <= "111";B <= "111";
					when 286=>
						R <= "111";G <= "111";B <= "111";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "111";G <= "111";B <= "111";
					when 289=>
						R <= "111";G <= "111";B <= "111";
					when 290=>
						R <= "101";G <= "100";B <= "011";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "110";
					when 296=>
						R <= "001";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "001";B <= "010";
					when 305=>
						R <= "110";G <= "111";B <= "111";
					when 306=>
						R <= "111";G <= "111";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "011";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "001";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "111";B <= "110";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "001";B <= "010";
					when 327=>
						R <= "110";G <= "111";B <= "111";
					when 328=>
						R <= "111";G <= "111";B <= "111";
					when 329=>
						R <= "100";G <= "011";B <= "010";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "011";G <= "100";B <= "100";
					when 340=>
						R <= "111";G <= "111";B <= "111";
					when 341=>
						R <= "111";G <= "111";B <= "111";
					when 342=>
						R <= "011";G <= "010";B <= "001";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "100";G <= "101";B <= "110";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "111";G <= "111";B <= "111";
					when 348=>
						R <= "111";G <= "111";B <= "111";
					when 349=>
						R <= "111";G <= "111";B <= "111";
					when 350=>
						R <= "111";G <= "111";B <= "111";
					when 351=>
						R <= "111";G <= "111";B <= "111";
					when 352=>
						R <= "111";G <= "111";B <= "111";
					when 353=>
						R <= "111";G <= "111";B <= "111";
					when 354=>
						R <= "111";G <= "111";B <= "111";
					when 355=>
						R <= "111";G <= "111";B <= "111";
					when 356=>
						R <= "001";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "011";G <= "100";B <= "101";
					when 363=>
						R <= "111";G <= "111";B <= "111";
					when 364=>
						R <= "111";G <= "111";B <= "111";
					when 365=>
						R <= "101";G <= "100";B <= "011";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "011";G <= "100";B <= "101";
					when 369=>
						R <= "111";G <= "111";B <= "111";
					when 370=>
						R <= "111";G <= "111";B <= "111";
					when 371=>
						R <= "101";G <= "100";B <= "011";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "011";G <= "100";B <= "100";
					when 375=>
						R <= "111";G <= "111";B <= "111";
					when 376=>
						R <= "111";G <= "111";B <= "111";
					when 377=>
						R <= "101";G <= "100";B <= "011";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 211=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "001";B <= "010";
					when 257=>
						R <= "111";G <= "111";B <= "111";
					when 258=>
						R <= "111";G <= "111";B <= "111";
					when 259=>
						R <= "011";G <= "010";B <= "001";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "011";G <= "100";B <= "100";
					when 268=>
						R <= "111";G <= "111";B <= "111";
					when 269=>
						R <= "111";G <= "110";B <= "110";
					when 270=>
						R <= "001";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "110";G <= "110";B <= "110";
					when 280=>
						R <= "111";G <= "111";B <= "111";
					when 281=>
						R <= "101";G <= "100";B <= "100";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "001";G <= "010";B <= "011";
					when 285=>
						R <= "111";G <= "111";B <= "111";
					when 286=>
						R <= "111";G <= "111";B <= "111";
					when 287=>
						R <= "111";G <= "111";B <= "111";
					when 288=>
						R <= "111";G <= "111";B <= "111";
					when 289=>
						R <= "111";G <= "111";B <= "111";
					when 290=>
						R <= "101";G <= "100";B <= "100";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "011";G <= "100";B <= "100";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "110";B <= "110";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "011";G <= "100";B <= "100";
					when 306=>
						R <= "111";G <= "111";B <= "111";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "101";G <= "100";B <= "100";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "011";G <= "100";B <= "100";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "111";G <= "110";B <= "110";
					when 316=>
						R <= "001";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "100";G <= "101";B <= "101";
					when 327=>
						R <= "111";G <= "111";B <= "111";
					when 328=>
						R <= "111";G <= "111";B <= "111";
					when 329=>
						R <= "001";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "001";
					when 340=>
						R <= "111";G <= "111";B <= "111";
					when 341=>
						R <= "111";G <= "111";B <= "111";
					when 342=>
						R <= "101";G <= "100";B <= "100";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "100";G <= "101";B <= "110";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "111";G <= "111";B <= "111";
					when 348=>
						R <= "111";G <= "111";B <= "111";
					when 349=>
						R <= "111";G <= "111";B <= "111";
					when 350=>
						R <= "111";G <= "111";B <= "111";
					when 351=>
						R <= "111";G <= "111";B <= "111";
					when 352=>
						R <= "111";G <= "111";B <= "111";
					when 353=>
						R <= "111";G <= "110";B <= "110";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "001";B <= "010";
					when 363=>
						R <= "111";G <= "111";B <= "111";
					when 364=>
						R <= "111";G <= "111";B <= "111";
					when 365=>
						R <= "011";G <= "010";B <= "001";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "001";B <= "010";
					when 369=>
						R <= "111";G <= "111";B <= "111";
					when 370=>
						R <= "111";G <= "111";B <= "111";
					when 371=>
						R <= "011";G <= "010";B <= "001";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "001";G <= "001";B <= "010";
					when 375=>
						R <= "111";G <= "111";B <= "111";
					when 376=>
						R <= "111";G <= "111";B <= "111";
					when 377=>
						R <= "011";G <= "010";B <= "001";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 212=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 213=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 214=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 215=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 216=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 217=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 218=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 219=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 220=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 221=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 222=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 223=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 224=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 225=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 226=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 227=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 228=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 229=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 230=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 231=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 232=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 233=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 234=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 235=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 236=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 237=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 238=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 239=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 240=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 241=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 242=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 243=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 244=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 245=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 246=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 247=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 248=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 249=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 250=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 251=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 252=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 253=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 254=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 255=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 256=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 257=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 258=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 259=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 260=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 261=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 262=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 263=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 264=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 265=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 266=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 267=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 268=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 269=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 270=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 271=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 272=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 273=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 274=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 275=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 276=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "010";G <= "010";B <= "010";
					when 310=>
						R <= "011";G <= "011";B <= "011";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "010";G <= "010";B <= "010";
					when 317=>
						R <= "100";G <= "100";B <= "100";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "011";G <= "011";B <= "010";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "101";G <= "110";B <= "110";
					when 327=>
						R <= "111";G <= "111";B <= "111";
					when 328=>
						R <= "111";G <= "111";B <= "111";
					when 329=>
						R <= "111";G <= "111";B <= "111";
					when 330=>
						R <= "011";G <= "011";B <= "010";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "001";G <= "001";B <= "001";
					when 335=>
						R <= "100";G <= "100";B <= "100";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "010";G <= "010";B <= "010";
					when 339=>
						R <= "011";G <= "011";B <= "011";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "011";G <= "011";B <= "010";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "100";G <= "101";B <= "101";
					when 364=>
						R <= "111";G <= "111";B <= "111";
					when 365=>
						R <= "111";G <= "111";B <= "111";
					when 366=>
						R <= "010";G <= "010";B <= "001";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "001";G <= "001";B <= "001";
					when 370=>
						R <= "111";G <= "111";B <= "110";
					when 371=>
						R <= "001";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "001";G <= "001";B <= "001";
					when 375=>
						R <= "111";G <= "111";B <= "111";
					when 376=>
						R <= "001";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 277=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "010";G <= "010";B <= "010";
					when 317=>
						R <= "100";G <= "101";B <= "101";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "101";G <= "101";B <= "100";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "101";G <= "110";B <= "110";
					when 326=>
						R <= "010";G <= "010";B <= "010";
					when 327=>
						R <= "001";G <= "001";B <= "001";
					when 328=>
						R <= "100";G <= "100";B <= "100";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "101";G <= "101";B <= "100";
					when 331=>
						R <= "010";G <= "010";B <= "001";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "001";G <= "001";B <= "001";
					when 335=>
						R <= "100";G <= "100";B <= "100";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "101";G <= "101";B <= "100";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "101";G <= "110";B <= "110";
					when 364=>
						R <= "000";G <= "000";B <= "001";
					when 365=>
						R <= "100";G <= "011";B <= "011";
					when 366=>
						R <= "011";G <= "011";B <= "010";
					when 367=>
						R <= "100";G <= "011";B <= "011";
					when 368=>
						R <= "010";G <= "010";B <= "010";
					when 369=>
						R <= "001";G <= "001";B <= "001";
					when 370=>
						R <= "110";G <= "110";B <= "101";
					when 371=>
						R <= "101";G <= "100";B <= "100";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "100";G <= "101";B <= "101";
					when 375=>
						R <= "101";G <= "101";B <= "101";
					when 376=>
						R <= "001";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 278=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "001";G <= "001";B <= "010";
					when 289=>
						R <= "111";G <= "111";B <= "111";
					when 290=>
						R <= "111";G <= "111";B <= "111";
					when 291=>
						R <= "110";G <= "110";B <= "110";
					when 292=>
						R <= "010";G <= "010";B <= "010";
					when 293=>
						R <= "111";G <= "111";B <= "111";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "111";B <= "111";
					when 296=>
						R <= "011";G <= "011";B <= "011";
					when 297=>
						R <= "010";G <= "010";B <= "010";
					when 298=>
						R <= "111";G <= "111";B <= "111";
					when 299=>
						R <= "111";G <= "111";B <= "111";
					when 300=>
						R <= "111";G <= "111";B <= "111";
					when 301=>
						R <= "101";G <= "100";B <= "100";
					when 302=>
						R <= "110";G <= "110";B <= "110";
					when 303=>
						R <= "010";G <= "010";B <= "010";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "101";G <= "110";B <= "110";
					when 306=>
						R <= "011";G <= "011";B <= "011";
					when 307=>
						R <= "111";G <= "111";B <= "111";
					when 308=>
						R <= "110";G <= "111";B <= "111";
					when 309=>
						R <= "010";G <= "011";B <= "011";
					when 310=>
						R <= "100";G <= "101";B <= "100";
					when 311=>
						R <= "010";G <= "010";B <= "010";
					when 312=>
						R <= "111";G <= "111";B <= "111";
					when 313=>
						R <= "111";G <= "111";B <= "111";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "100";G <= "100";B <= "100";
					when 316=>
						R <= "010";G <= "010";B <= "011";
					when 317=>
						R <= "111";G <= "111";B <= "111";
					when 318=>
						R <= "111";G <= "111";B <= "111";
					when 319=>
						R <= "111";G <= "111";B <= "111";
					when 320=>
						R <= "010";G <= "010";B <= "010";
					when 321=>
						R <= "101";G <= "101";B <= "101";
					when 322=>
						R <= "111";G <= "111";B <= "111";
					when 323=>
						R <= "110";G <= "110";B <= "101";
					when 324=>
						R <= "001";G <= "001";B <= "001";
					when 325=>
						R <= "100";G <= "100";B <= "100";
					when 326=>
						R <= "010";G <= "010";B <= "010";
					when 327=>
						R <= "110";G <= "110";B <= "111";
					when 328=>
						R <= "100";G <= "100";B <= "100";
					when 329=>
						R <= "100";G <= "100";B <= "100";
					when 330=>
						R <= "001";G <= "001";B <= "001";
					when 331=>
						R <= "100";G <= "100";B <= "100";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "001";G <= "001";B <= "001";
					when 335=>
						R <= "100";G <= "100";B <= "100";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "010";G <= "010";B <= "010";
					when 339=>
						R <= "100";G <= "101";B <= "100";
					when 340=>
						R <= "010";G <= "010";B <= "010";
					when 341=>
						R <= "011";G <= "011";B <= "011";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "011";G <= "100";B <= "100";
					when 344=>
						R <= "011";G <= "011";B <= "011";
					when 345=>
						R <= "101";G <= "101";B <= "100";
					when 346=>
						R <= "111";G <= "111";B <= "111";
					when 347=>
						R <= "110";G <= "110";B <= "101";
					when 348=>
						R <= "011";G <= "100";B <= "100";
					when 349=>
						R <= "111";G <= "111";B <= "111";
					when 350=>
						R <= "111";G <= "111";B <= "111";
					when 351=>
						R <= "010";G <= "010";B <= "010";
					when 352=>
						R <= "001";G <= "001";B <= "010";
					when 353=>
						R <= "111";G <= "111";B <= "111";
					when 354=>
						R <= "111";G <= "111";B <= "111";
					when 355=>
						R <= "111";G <= "111";B <= "111";
					when 356=>
						R <= "000";G <= "000";B <= "001";
					when 357=>
						R <= "010";G <= "010";B <= "010";
					when 358=>
						R <= "111";G <= "111";B <= "111";
					when 359=>
						R <= "111";G <= "111";B <= "111";
					when 360=>
						R <= "111";G <= "111";B <= "111";
					when 361=>
						R <= "010";G <= "010";B <= "010";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "001";B <= "010";
					when 364=>
						R <= "111";G <= "111";B <= "111";
					when 365=>
						R <= "100";G <= "100";B <= "100";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "011";G <= "011";B <= "011";
					when 368=>
						R <= "010";G <= "010";B <= "010";
					when 369=>
						R <= "001";G <= "001";B <= "001";
					when 370=>
						R <= "100";G <= "100";B <= "100";
					when 371=>
						R <= "101";G <= "110";B <= "101";
					when 372=>
						R <= "001";G <= "001";B <= "000";
					when 373=>
						R <= "001";G <= "001";B <= "001";
					when 374=>
						R <= "101";G <= "110";B <= "101";
					when 375=>
						R <= "110";G <= "110";B <= "110";
					when 376=>
						R <= "001";G <= "000";B <= "001";
					when 377=>
						R <= "010";G <= "001";B <= "001";
					when 378=>
						R <= "111";G <= "111";B <= "111";
					when 379=>
						R <= "111";G <= "111";B <= "111";
					when 380=>
						R <= "110";G <= "110";B <= "101";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 279=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "011";G <= "100";B <= "100";
					when 289=>
						R <= "001";G <= "010";B <= "010";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "100";G <= "101";B <= "101";
					when 293=>
						R <= "001";G <= "010";B <= "011";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "001";G <= "001";B <= "010";
					when 296=>
						R <= "101";G <= "101";B <= "110";
					when 297=>
						R <= "010";G <= "010";B <= "010";
					when 298=>
						R <= "101";G <= "100";B <= "100";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "001";G <= "000";B <= "000";
					when 301=>
						R <= "101";G <= "101";B <= "101";
					when 302=>
						R <= "001";G <= "001";B <= "001";
					when 303=>
						R <= "100";G <= "100";B <= "100";
					when 304=>
						R <= "001";G <= "001";B <= "001";
					when 305=>
						R <= "100";G <= "100";B <= "100";
					when 306=>
						R <= "010";G <= "010";B <= "010";
					when 307=>
						R <= "100";G <= "101";B <= "101";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "001";G <= "010";B <= "011";
					when 310=>
						R <= "100";G <= "101";B <= "101";
					when 311=>
						R <= "011";G <= "011";B <= "011";
					when 312=>
						R <= "010";G <= "010";B <= "010";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "010";G <= "010";B <= "001";
					when 315=>
						R <= "101";G <= "101";B <= "100";
					when 316=>
						R <= "010";G <= "010";B <= "010";
					when 317=>
						R <= "100";G <= "101";B <= "101";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "011";G <= "100";B <= "100";
					when 320=>
						R <= "011";G <= "011";B <= "011";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "101";G <= "101";B <= "100";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "010";G <= "010";B <= "010";
					when 325=>
						R <= "011";G <= "011";B <= "011";
					when 326=>
						R <= "100";G <= "100";B <= "101";
					when 327=>
						R <= "000";G <= "001";B <= "001";
					when 328=>
						R <= "001";G <= "001";B <= "001";
					when 329=>
						R <= "100";G <= "100";B <= "100";
					when 330=>
						R <= "001";G <= "001";B <= "001";
					when 331=>
						R <= "100";G <= "100";B <= "100";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "001";G <= "001";B <= "001";
					when 335=>
						R <= "100";G <= "100";B <= "100";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "010";G <= "010";B <= "010";
					when 339=>
						R <= "100";G <= "100";B <= "100";
					when 340=>
						R <= "010";G <= "010";B <= "010";
					when 341=>
						R <= "011";G <= "011";B <= "011";
					when 342=>
						R <= "000";G <= "000";B <= "001";
					when 343=>
						R <= "011";G <= "011";B <= "100";
					when 344=>
						R <= "011";G <= "011";B <= "011";
					when 345=>
						R <= "001";G <= "000";B <= "000";
					when 346=>
						R <= "101";G <= "101";B <= "100";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "001";G <= "010";B <= "011";
					when 349=>
						R <= "111";G <= "111";B <= "111";
					when 350=>
						R <= "001";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "100";G <= "101";B <= "101";
					when 353=>
						R <= "111";G <= "111";B <= "111";
					when 354=>
						R <= "111";G <= "111";B <= "111";
					when 355=>
						R <= "111";G <= "111";B <= "111";
					when 356=>
						R <= "010";G <= "010";B <= "010";
					when 357=>
						R <= "010";G <= "010";B <= "010";
					when 358=>
						R <= "101";G <= "100";B <= "100";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "100";G <= "011";B <= "011";
					when 361=>
						R <= "011";G <= "011";B <= "011";
					when 362=>
						R <= "010";G <= "010";B <= "010";
					when 363=>
						R <= "110";G <= "111";B <= "111";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "011";G <= "011";B <= "011";
					when 366=>
						R <= "011";G <= "011";B <= "011";
					when 367=>
						R <= "101";G <= "101";B <= "101";
					when 368=>
						R <= "000";G <= "000";B <= "001";
					when 369=>
						R <= "001";G <= "001";B <= "001";
					when 370=>
						R <= "100";G <= "100";B <= "100";
					when 371=>
						R <= "010";G <= "010";B <= "001";
					when 372=>
						R <= "011";G <= "011";B <= "011";
					when 373=>
						R <= "011";G <= "011";B <= "011";
					when 374=>
						R <= "010";G <= "010";B <= "010";
					when 375=>
						R <= "101";G <= "101";B <= "101";
					when 376=>
						R <= "001";G <= "000";B <= "001";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "011";G <= "011";B <= "100";
					when 379=>
						R <= "111";G <= "111";B <= "111";
					when 380=>
						R <= "111";G <= "110";B <= "101";
					when 381=>
						R <= "001";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 280=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "011";G <= "100";B <= "100";
					when 289=>
						R <= "011";G <= "011";B <= "011";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "011";G <= "100";B <= "100";
					when 293=>
						R <= "011";G <= "011";B <= "100";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "001";G <= "001";B <= "010";
					when 296=>
						R <= "101";G <= "101";B <= "110";
					when 297=>
						R <= "010";G <= "010";B <= "010";
					when 298=>
						R <= "101";G <= "100";B <= "100";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "010";G <= "001";B <= "000";
					when 301=>
						R <= "110";G <= "101";B <= "101";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "101";G <= "101";B <= "101";
					when 304=>
						R <= "101";G <= "101";B <= "101";
					when 305=>
						R <= "010";G <= "010";B <= "001";
					when 306=>
						R <= "010";G <= "010";B <= "010";
					when 307=>
						R <= "100";G <= "101";B <= "101";
					when 308=>
						R <= "000";G <= "000";B <= "001";
					when 309=>
						R <= "001";G <= "010";B <= "011";
					when 310=>
						R <= "100";G <= "100";B <= "101";
					when 311=>
						R <= "100";G <= "011";B <= "011";
					when 312=>
						R <= "010";G <= "010";B <= "001";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "010";G <= "010";B <= "001";
					when 315=>
						R <= "101";G <= "100";B <= "100";
					when 316=>
						R <= "010";G <= "010";B <= "010";
					when 317=>
						R <= "100";G <= "101";B <= "101";
					when 318=>
						R <= "000";G <= "000";B <= "001";
					when 319=>
						R <= "011";G <= "100";B <= "100";
					when 320=>
						R <= "011";G <= "011";B <= "011";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "101";G <= "101";B <= "100";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "001";G <= "001";B <= "001";
					when 325=>
						R <= "100";G <= "100";B <= "100";
					when 326=>
						R <= "011";G <= "100";B <= "100";
					when 327=>
						R <= "011";G <= "011";B <= "011";
					when 328=>
						R <= "101";G <= "101";B <= "100";
					when 329=>
						R <= "101";G <= "101";B <= "100";
					when 330=>
						R <= "100";G <= "011";B <= "011";
					when 331=>
						R <= "010";G <= "010";B <= "010";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "001";B <= "001";
					when 335=>
						R <= "100";G <= "100";B <= "101";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "010";G <= "010";B <= "010";
					when 339=>
						R <= "100";G <= "100";B <= "101";
					when 340=>
						R <= "010";G <= "010";B <= "010";
					when 341=>
						R <= "011";G <= "011";B <= "100";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "011";G <= "100";B <= "100";
					when 344=>
						R <= "100";G <= "011";B <= "011";
					when 345=>
						R <= "001";G <= "000";B <= "000";
					when 346=>
						R <= "101";G <= "101";B <= "100";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "001";
					when 349=>
						R <= "000";G <= "000";B <= "001";
					when 350=>
						R <= "111";G <= "111";B <= "110";
					when 351=>
						R <= "100";G <= "011";B <= "010";
					when 352=>
						R <= "011";G <= "100";B <= "100";
					when 353=>
						R <= "010";G <= "010";B <= "010";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "010";G <= "010";B <= "011";
					when 358=>
						R <= "101";G <= "100";B <= "100";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "100";G <= "011";B <= "011";
					when 361=>
						R <= "011";G <= "011";B <= "011";
					when 362=>
						R <= "011";G <= "100";B <= "100";
					when 363=>
						R <= "011";G <= "011";B <= "100";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "101";G <= "101";B <= "101";
					when 367=>
						R <= "011";G <= "011";B <= "011";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "001";G <= "001";B <= "010";
					when 370=>
						R <= "100";G <= "100";B <= "100";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "110";G <= "110";B <= "101";
					when 373=>
						R <= "110";G <= "110";B <= "110";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "101";G <= "110";B <= "110";
					when 376=>
						R <= "001";G <= "000";B <= "001";
					when 377=>
						R <= "101";G <= "100";B <= "101";
					when 378=>
						R <= "101";G <= "100";B <= "101";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "110";G <= "110";B <= "101";
					when 381=>
						R <= "001";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 281=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "111";G <= "111";B <= "111";
					when 290=>
						R <= "111";G <= "111";B <= "111";
					when 291=>
						R <= "110";G <= "110";B <= "101";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "110";G <= "111";B <= "111";
					when 294=>
						R <= "111";G <= "111";B <= "111";
					when 295=>
						R <= "111";G <= "111";B <= "111";
					when 296=>
						R <= "000";G <= "001";B <= "001";
					when 297=>
						R <= "010";G <= "010";B <= "010";
					when 298=>
						R <= "111";G <= "111";B <= "111";
					when 299=>
						R <= "111";G <= "111";B <= "111";
					when 300=>
						R <= "111";G <= "111";B <= "111";
					when 301=>
						R <= "010";G <= "010";B <= "010";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "011";G <= "011";B <= "100";
					when 304=>
						R <= "110";G <= "110";B <= "101";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "010";G <= "010";B <= "010";
					when 307=>
						R <= "100";G <= "101";B <= "101";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "001";G <= "010";B <= "011";
					when 310=>
						R <= "100";G <= "101";B <= "101";
					when 311=>
						R <= "001";G <= "001";B <= "001";
					when 312=>
						R <= "111";G <= "111";B <= "111";
					when 313=>
						R <= "111";G <= "111";B <= "111";
					when 314=>
						R <= "111";G <= "111";B <= "111";
					when 315=>
						R <= "101";G <= "101";B <= "100";
					when 316=>
						R <= "010";G <= "010";B <= "010";
					when 317=>
						R <= "100";G <= "100";B <= "101";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "011";G <= "100";B <= "100";
					when 320=>
						R <= "011";G <= "011";B <= "011";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "111";G <= "111";B <= "110";
					when 323=>
						R <= "110";G <= "111";B <= "110";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "100";G <= "101";B <= "101";
					when 326=>
						R <= "010";G <= "010";B <= "010";
					when 327=>
						R <= "101";G <= "101";B <= "101";
					when 328=>
						R <= "011";G <= "011";B <= "011";
					when 329=>
						R <= "100";G <= "011";B <= "011";
					when 330=>
						R <= "101";G <= "100";B <= "100";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "001";G <= "001";B <= "010";
					when 335=>
						R <= "111";G <= "111";B <= "111";
					when 336=>
						R <= "111";G <= "111";B <= "111";
					when 337=>
						R <= "111";G <= "111";B <= "111";
					when 338=>
						R <= "011";G <= "011";B <= "011";
					when 339=>
						R <= "100";G <= "101";B <= "101";
					when 340=>
						R <= "001";G <= "001";B <= "010";
					when 341=>
						R <= "111";G <= "111";B <= "111";
					when 342=>
						R <= "111";G <= "111";B <= "111";
					when 343=>
						R <= "111";G <= "111";B <= "111";
					when 344=>
						R <= "011";G <= "011";B <= "011";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "111";G <= "111";B <= "110";
					when 347=>
						R <= "110";G <= "111";B <= "110";
					when 348=>
						R <= "011";G <= "100";B <= "101";
					when 349=>
						R <= "111";G <= "111";B <= "111";
					when 350=>
						R <= "111";G <= "111";B <= "111";
					when 351=>
						R <= "010";G <= "010";B <= "001";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "111";G <= "111";B <= "111";
					when 354=>
						R <= "111";G <= "111";B <= "111";
					when 355=>
						R <= "111";G <= "110";B <= "110";
					when 356=>
						R <= "000";G <= "000";B <= "001";
					when 357=>
						R <= "010";G <= "010";B <= "010";
					when 358=>
						R <= "101";G <= "100";B <= "100";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "100";G <= "011";B <= "011";
					when 361=>
						R <= "011";G <= "011";B <= "011";
					when 362=>
						R <= "001";G <= "001";B <= "001";
					when 363=>
						R <= "111";G <= "111";B <= "111";
					when 364=>
						R <= "111";G <= "111";B <= "111";
					when 365=>
						R <= "111";G <= "111";B <= "111";
					when 366=>
						R <= "011";G <= "011";B <= "011";
					when 367=>
						R <= "111";G <= "111";B <= "111";
					when 368=>
						R <= "110";G <= "110";B <= "111";
					when 369=>
						R <= "010";G <= "010";B <= "010";
					when 370=>
						R <= "100";G <= "100";B <= "100";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "011";G <= "100";B <= "011";
					when 373=>
						R <= "011";G <= "011";B <= "011";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "101";G <= "101";B <= "110";
					when 376=>
						R <= "001";G <= "000";B <= "001";
					when 377=>
						R <= "100";G <= "011";B <= "100";
					when 378=>
						R <= "111";G <= "111";B <= "111";
					when 379=>
						R <= "111";G <= "111";B <= "111";
					when 380=>
						R <= "111";G <= "110";B <= "101";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 282=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "001";
					when 297=>
						R <= "001";G <= "010";B <= "011";
					when 298=>
						R <= "101";G <= "100";B <= "100";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "011";G <= "100";B <= "100";
					when 304=>
						R <= "011";G <= "011";B <= "010";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "100";G <= "100";B <= "011";
					when 315=>
						R <= "011";G <= "011";B <= "010";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "101";G <= "110";B <= "110";
					when 327=>
						R <= "111";G <= "111";B <= "111";
					when 328=>
						R <= "111";G <= "111";B <= "111";
					when 329=>
						R <= "111";G <= "110";B <= "110";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 283=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "001";G <= "010";B <= "011";
					when 298=>
						R <= "101";G <= "100";B <= "100";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "101";G <= "110";B <= "110";
					when 303=>
						R <= "110";G <= "111";B <= "111";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "010";G <= "010";B <= "010";
					when 312=>
						R <= "111";G <= "111";B <= "111";
					when 313=>
						R <= "111";G <= "111";B <= "111";
					when 314=>
						R <= "111";G <= "110";B <= "110";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 284=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 285=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 286=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 287=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 288=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 289=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 290=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 291=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 292=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 293=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 294=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 295=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 296=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 297=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 298=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when 299=>
				case col is 
					when 240=>
						R <= "000";G <= "000";B <= "000";
					when 241=>
						R <= "000";G <= "000";B <= "000";
					when 242=>
						R <= "000";G <= "000";B <= "000";
					when 243=>
						R <= "000";G <= "000";B <= "000";
					when 244=>
						R <= "000";G <= "000";B <= "000";
					when 245=>
						R <= "000";G <= "000";B <= "000";
					when 246=>
						R <= "000";G <= "000";B <= "000";
					when 247=>
						R <= "000";G <= "000";B <= "000";
					when 248=>
						R <= "000";G <= "000";B <= "000";
					when 249=>
						R <= "000";G <= "000";B <= "000";
					when 250=>
						R <= "000";G <= "000";B <= "000";
					when 251=>
						R <= "000";G <= "000";B <= "000";
					when 252=>
						R <= "000";G <= "000";B <= "000";
					when 253=>
						R <= "000";G <= "000";B <= "000";
					when 254=>
						R <= "000";G <= "000";B <= "000";
					when 255=>
						R <= "000";G <= "000";B <= "000";
					when 256=>
						R <= "000";G <= "000";B <= "000";
					when 257=>
						R <= "000";G <= "000";B <= "000";
					when 258=>
						R <= "000";G <= "000";B <= "000";
					when 259=>
						R <= "000";G <= "000";B <= "000";
					when 260=>
						R <= "000";G <= "000";B <= "000";
					when 261=>
						R <= "000";G <= "000";B <= "000";
					when 262=>
						R <= "000";G <= "000";B <= "000";
					when 263=>
						R <= "000";G <= "000";B <= "000";
					when 264=>
						R <= "000";G <= "000";B <= "000";
					when 265=>
						R <= "000";G <= "000";B <= "000";
					when 266=>
						R <= "000";G <= "000";B <= "000";
					when 267=>
						R <= "000";G <= "000";B <= "000";
					when 268=>
						R <= "000";G <= "000";B <= "000";
					when 269=>
						R <= "000";G <= "000";B <= "000";
					when 270=>
						R <= "000";G <= "000";B <= "000";
					when 271=>
						R <= "000";G <= "000";B <= "000";
					when 272=>
						R <= "000";G <= "000";B <= "000";
					when 273=>
						R <= "000";G <= "000";B <= "000";
					when 274=>
						R <= "000";G <= "000";B <= "000";
					when 275=>
						R <= "000";G <= "000";B <= "000";
					when 276=>
						R <= "000";G <= "000";B <= "000";
					when 277=>
						R <= "000";G <= "000";B <= "000";
					when 278=>
						R <= "000";G <= "000";B <= "000";
					when 279=>
						R <= "000";G <= "000";B <= "000";
					when 280=>
						R <= "000";G <= "000";B <= "000";
					when 281=>
						R <= "000";G <= "000";B <= "000";
					when 282=>
						R <= "000";G <= "000";B <= "000";
					when 283=>
						R <= "000";G <= "000";B <= "000";
					when 284=>
						R <= "000";G <= "000";B <= "000";
					when 285=>
						R <= "000";G <= "000";B <= "000";
					when 286=>
						R <= "000";G <= "000";B <= "000";
					when 287=>
						R <= "000";G <= "000";B <= "000";
					when 288=>
						R <= "000";G <= "000";B <= "000";
					when 289=>
						R <= "000";G <= "000";B <= "000";
					when 290=>
						R <= "000";G <= "000";B <= "000";
					when 291=>
						R <= "000";G <= "000";B <= "000";
					when 292=>
						R <= "000";G <= "000";B <= "000";
					when 293=>
						R <= "000";G <= "000";B <= "000";
					when 294=>
						R <= "000";G <= "000";B <= "000";
					when 295=>
						R <= "000";G <= "000";B <= "000";
					when 296=>
						R <= "000";G <= "000";B <= "000";
					when 297=>
						R <= "000";G <= "000";B <= "000";
					when 298=>
						R <= "000";G <= "000";B <= "000";
					when 299=>
						R <= "000";G <= "000";B <= "000";
					when 300=>
						R <= "000";G <= "000";B <= "000";
					when 301=>
						R <= "000";G <= "000";B <= "000";
					when 302=>
						R <= "000";G <= "000";B <= "000";
					when 303=>
						R <= "000";G <= "000";B <= "000";
					when 304=>
						R <= "000";G <= "000";B <= "000";
					when 305=>
						R <= "000";G <= "000";B <= "000";
					when 306=>
						R <= "000";G <= "000";B <= "000";
					when 307=>
						R <= "000";G <= "000";B <= "000";
					when 308=>
						R <= "000";G <= "000";B <= "000";
					when 309=>
						R <= "000";G <= "000";B <= "000";
					when 310=>
						R <= "000";G <= "000";B <= "000";
					when 311=>
						R <= "000";G <= "000";B <= "000";
					when 312=>
						R <= "000";G <= "000";B <= "000";
					when 313=>
						R <= "000";G <= "000";B <= "000";
					when 314=>
						R <= "000";G <= "000";B <= "000";
					when 315=>
						R <= "000";G <= "000";B <= "000";
					when 316=>
						R <= "000";G <= "000";B <= "000";
					when 317=>
						R <= "000";G <= "000";B <= "000";
					when 318=>
						R <= "000";G <= "000";B <= "000";
					when 319=>
						R <= "000";G <= "000";B <= "000";
					when 320=>
						R <= "000";G <= "000";B <= "000";
					when 321=>
						R <= "000";G <= "000";B <= "000";
					when 322=>
						R <= "000";G <= "000";B <= "000";
					when 323=>
						R <= "000";G <= "000";B <= "000";
					when 324=>
						R <= "000";G <= "000";B <= "000";
					when 325=>
						R <= "000";G <= "000";B <= "000";
					when 326=>
						R <= "000";G <= "000";B <= "000";
					when 327=>
						R <= "000";G <= "000";B <= "000";
					when 328=>
						R <= "000";G <= "000";B <= "000";
					when 329=>
						R <= "000";G <= "000";B <= "000";
					when 330=>
						R <= "000";G <= "000";B <= "000";
					when 331=>
						R <= "000";G <= "000";B <= "000";
					when 332=>
						R <= "000";G <= "000";B <= "000";
					when 333=>
						R <= "000";G <= "000";B <= "000";
					when 334=>
						R <= "000";G <= "000";B <= "000";
					when 335=>
						R <= "000";G <= "000";B <= "000";
					when 336=>
						R <= "000";G <= "000";B <= "000";
					when 337=>
						R <= "000";G <= "000";B <= "000";
					when 338=>
						R <= "000";G <= "000";B <= "000";
					when 339=>
						R <= "000";G <= "000";B <= "000";
					when 340=>
						R <= "000";G <= "000";B <= "000";
					when 341=>
						R <= "000";G <= "000";B <= "000";
					when 342=>
						R <= "000";G <= "000";B <= "000";
					when 343=>
						R <= "000";G <= "000";B <= "000";
					when 344=>
						R <= "000";G <= "000";B <= "000";
					when 345=>
						R <= "000";G <= "000";B <= "000";
					when 346=>
						R <= "000";G <= "000";B <= "000";
					when 347=>
						R <= "000";G <= "000";B <= "000";
					when 348=>
						R <= "000";G <= "000";B <= "000";
					when 349=>
						R <= "000";G <= "000";B <= "000";
					when 350=>
						R <= "000";G <= "000";B <= "000";
					when 351=>
						R <= "000";G <= "000";B <= "000";
					when 352=>
						R <= "000";G <= "000";B <= "000";
					when 353=>
						R <= "000";G <= "000";B <= "000";
					when 354=>
						R <= "000";G <= "000";B <= "000";
					when 355=>
						R <= "000";G <= "000";B <= "000";
					when 356=>
						R <= "000";G <= "000";B <= "000";
					when 357=>
						R <= "000";G <= "000";B <= "000";
					when 358=>
						R <= "000";G <= "000";B <= "000";
					when 359=>
						R <= "000";G <= "000";B <= "000";
					when 360=>
						R <= "000";G <= "000";B <= "000";
					when 361=>
						R <= "000";G <= "000";B <= "000";
					when 362=>
						R <= "000";G <= "000";B <= "000";
					when 363=>
						R <= "000";G <= "000";B <= "000";
					when 364=>
						R <= "000";G <= "000";B <= "000";
					when 365=>
						R <= "000";G <= "000";B <= "000";
					when 366=>
						R <= "000";G <= "000";B <= "000";
					when 367=>
						R <= "000";G <= "000";B <= "000";
					when 368=>
						R <= "000";G <= "000";B <= "000";
					when 369=>
						R <= "000";G <= "000";B <= "000";
					when 370=>
						R <= "000";G <= "000";B <= "000";
					when 371=>
						R <= "000";G <= "000";B <= "000";
					when 372=>
						R <= "000";G <= "000";B <= "000";
					when 373=>
						R <= "000";G <= "000";B <= "000";
					when 374=>
						R <= "000";G <= "000";B <= "000";
					when 375=>
						R <= "000";G <= "000";B <= "000";
					when 376=>
						R <= "000";G <= "000";B <= "000";
					when 377=>
						R <= "000";G <= "000";B <= "000";
					when 378=>
						R <= "000";G <= "000";B <= "000";
					when 379=>
						R <= "000";G <= "000";B <= "000";
					when 380=>
						R <= "000";G <= "000";B <= "000";
					when 381=>
						R <= "000";G <= "000";B <= "000";
					when 382=>
						R <= "000";G <= "000";B <= "000";
					when 383=>
						R <= "000";G <= "000";B <= "000";
					when 384=>
						R <= "000";G <= "000";B <= "000";
					when 385=>
						R <= "000";G <= "000";B <= "000";
					when 386=>
						R <= "000";G <= "000";B <= "000";
					when 387=>
						R <= "000";G <= "000";B <= "000";
					when 388=>
						R <= "000";G <= "000";B <= "000";
					when 389=>
						R <= "000";G <= "000";B <= "000";
					when 390=>
						R <= "000";G <= "000";B <= "000";
					when 391=>
						R <= "000";G <= "000";B <= "000";
					when 392=>
						R <= "000";G <= "000";B <= "000";
					when 393=>
						R <= "000";G <= "000";B <= "000";
					when 394=>
						R <= "000";G <= "000";B <= "000";
					when 395=>
						R <= "000";G <= "000";B <= "000";
					when 396=>
						R <= "000";G <= "000";B <= "000";
					when 397=>
						R <= "000";G <= "000";B <= "000";
					when 398=>
						R <= "000";G <= "000";B <= "000";
					when 399=>
						R <= "000";G <= "000";B <= "000";
					when others=>
						R <= "000";G <= "000";B <= "000";		
				end case;
			when others=>
				R<="000";G<="000";B<="000";
		end case;

		if col>=656 and col<=752 then
			Hs<='0';
		else
			Hs<='1';
		end if;
		if row>=490 and row<=491 then
			Vs<='0';
		else
			Vs<='1';
		end if;
		if col=799 then
			col:=0;
			if row=524 then
				row:=0;
			else
				row:=row+1;
			end if;
		else
			col:=col+1;
		end if;
	end if;
end process;

end Behavioral;